// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_RAL_ST_MACROS_SV__
`define __UVME_RAL_ST_MACROS_SV__





`endif // __UVME_RAL_ST_MACROS_SV__
