// Copyright 2021 OpenHW Group
// Copyright 2021 Datum Technology Corporation
// Copyright 2021 Silicon Labs
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVML_RAL_TDEFS_SV__
`define __UVML_RAL_TDEFS_SV__


/**
 *
 */
typedef enum {
    UVML_RAL_MEM_DEFAULT_VAL_X     , ///<
    UVML_RAL_MEM_DEFAULT_VAL_0     , ///<
    UVML_RAL_MEM_DEFAULT_VAL_CONST , ///<
    UVML_RAL_MEM_DEFAULT_VAL_INCR  , ///<
    UVML_RAL_MEM_DEFAULT_VAL_RANDOM  ///<
} uvml_ral_mem_default_val_enum;


`endif // __UVML_RAL_TDEFS_SV__
