// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVML_RAL_CONSTANTS_SV__
`define __UVML_RAL_CONSTANTS_SV__





`endif // __UVML_RAL_CONSTANTS_SV__
